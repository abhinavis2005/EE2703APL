.circuit
R1   1                                  GND     1
.end
